module nor_gate(output o2,input a2,b2);
nor nor_gate(o2,a2,b2);
endmodule