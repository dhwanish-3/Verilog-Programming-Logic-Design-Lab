module nor_1(output o,input a);
nor g1(o,a);
endmodule