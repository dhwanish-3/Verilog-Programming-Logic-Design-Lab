module array_nor_gate(output [0:15]o,input [0:15]a,b);
nor g1(o[0],a[0],b[0]);
nor g2(o[1],a[1],b[1]);
nor g3(o[2],a[2],b[2]);
nor g4(o[3],a[3],b[3]);
nor g5(o[4],a[4],b[4]);
nor g6(o[5],a[5],b[5]);
nor g7(o[6],a[6],b[6]);
nor g8(o[7],a[7],b[7]);
nor g9(o[8],a[8],b[8]);
nor gq(o[9],a[9],b[9]);
nor gw(o[10],a[10],b[10]);
nor ge(o[11],a[11],b[11]);
nor gr(o[12],a[12],b[12]);
nor gy(o[13],a[13],b[13]);
nor gt(o[14],a[14],b[14]);
nor gu(o[15],a[15],b[15]);
endmodule
