module inverter_data(o1,i1);
output o1;
input i1;
assign o1=~i1;
endmodule
