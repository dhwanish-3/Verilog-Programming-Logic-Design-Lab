module clockDLatch_A(input d,pre,clr,output q,qbar);

endmodule
