module nand_1(output o,input a);
nand g1(o,a);
endmodule