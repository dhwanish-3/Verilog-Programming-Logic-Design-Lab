module array_not_data(output [0:15]o,input [0:15]a);
not g1(o[0],a[0]);
not g2(o[1],a[1]);
not g3(o[2],a[2]);
not g4(o[3],a[3]);
not g5(o[4],a[4]);
not g6(o[5],a[5]);
not g7(o[6],a[6]);
not g8(o[7],a[7]);
not g9(o[8],a[8]);
not gq(o[9],a[9]);
not gw(o[10],a[10]);
not ge(o[11],a[11]);
not gr(o[12],a[12]);
not gy(o[13],a[13]);
not gt(o[14],a[14]);
not gu(o[15],a[15]);
endmodule
