module inverter_gate(output o1,input i1);
not inverter_gate(o1,i1);
endmodule
