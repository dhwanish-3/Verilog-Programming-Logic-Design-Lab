module array_and(output [0:15]o,input [0:15]a,b);
assign o=a&b;
endmodule
