module nand_not_data(output o,input a);
assign o=~a;
endmodule
